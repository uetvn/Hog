--------------------------------------------------------------------------------
-- Project name   : Human detection by HOG
-- File name      : hog_block_8x8.vhd
-- Created date   : Mon 24 Apr 2017
-- Author         : Huy Hung Ho
-- Last modified  : Mon 24 Apr 2017
-- Desc           :
--------------------------------------------------------------------------------
package X is
    function 




library IEEE;
use IEEE.std_logic_1164.all;

entity hog_block_8x8 is
	Port (
        
	);
end hog_block_8x8;

architecture behav of hog_block_8x8 is

begin

end behav;

