--------------------------------------------------------------------------------
-- Project name   : Human detection by HOG
-- File name      : src/lut.vhd
-- Created date   : Monday 07/03/17
-- Author         : Huy Hung Ho
-- Last modified  : Monday 07/03/17
-- Desc           :
--------------------------------------------------------------------------------

Library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.math_real.all;
library std;
use std.textio.all;

Entity lut_16x16 is
    port(
            clk:        IN std_logic;
            enable:     IN std_logic;
            dx:         IN real;
            dy:         IN real;
            magnit:     OUT real;
            angle:      OUT real
	);
End lut_16x16;

Architecture Behavioral of lut_16x16 is
    Constant mem_depth: integer := 2 * 16 * 16;
    Type     RAM is array (integer range <>) of real range 0.0 to 256.0;
    Signal   mem: RAM(0 to mem_depth - 1)
        := (1.4142,2.2361,3.1623,4.1231,5.099,6.0828,7.0711,8.0623,9.0554,10.05,11.045,12.042,13.038,14.036,15.033,16.031,
2.2361,2.8284,3.6056,4.4721,5.3852,6.3246,7.2801,8.2462,9.2195,10.198,11.18,12.166,13.153,14.142,15.133,16.125,
3.1623,3.6056,4.2426,5.0,5.831,6.7082,7.6158,8.544,9.4868,10.44,11.402,12.369,13.342,14.318,15.297,16.279,
4.1231,4.4721,5.0,5.6569,6.4031,7.2111,8.0623,8.9443,9.8489,10.77,11.705,12.649,13.601,14.56,15.524,16.492,
5.099,5.3852,5.831,6.4031,7.0711,7.8102,8.6023,9.434,10.296,11.18,12.083,13.0,13.928,14.866,15.811,16.763,
6.0828,6.3246,6.7082,7.2111,7.8102,8.4853,9.2195,10.0,10.817,11.662,12.53,13.416,14.318,15.232,16.155,17.088,
7.0711,7.2801,7.6158,8.0623,8.6023,9.2195,9.8995,10.63,11.402,12.207,13.038,13.892,14.765,15.652,16.553,17.464,
8.0623,8.2462,8.544,8.9443,9.434,10.0,10.63,11.314,12.042,12.806,13.601,14.422,15.264,16.125,17.0,17.889,
9.0554,9.2195,9.4868,9.8489,10.296,10.817,11.402,12.042,12.728,13.454,14.213,15.0,15.811,16.643,17.493,18.358,
10.05,10.198,10.44,10.77,11.18,11.662,12.207,12.806,13.454,14.142,14.866,15.62,16.401,17.205,18.028,18.868,
11.045,11.18,11.402,11.705,12.083,12.53,13.038,13.601,14.213,14.866,15.556,16.279,17.029,17.804,18.601,19.416,
12.042,12.166,12.369,12.649,13.0,13.416,13.892,14.422,15.0,15.62,16.279,16.971,17.692,18.439,19.209,20.0,
13.038,13.153,13.342,13.601,13.928,14.318,14.765,15.264,15.811,16.401,17.029,17.692,18.385,19.105,19.849,20.616,
14.036,14.142,14.318,14.56,14.866,15.232,15.652,16.125,16.643,17.205,17.804,18.439,19.105,19.799,20.518,21.26,
15.033,15.133,15.297,15.524,15.811,16.155,16.553,17.0,17.493,18.028,18.601,19.209,19.849,20.518,21.213,21.932,
16.031,16.125,16.279,16.492,16.763,17.088,17.464,17.889,18.358,18.868,19.416,20.0,20.616,21.26,21.932,22.627,
			0.7854, 0.4636, 0.3218, 0.2450, 0.1974, 0.1651, 0.1419, 0.1244, 0.1107, 0.0997, 0.0907, 0.0831, 0.0768, 0.0713, 0.0666, 0.0624, 1.1072,
0.7854, 0.5880, 0.4636, 0.3805, 0.3218, 0.2783, 0.2450, 0.2187, 0.1974, 0.1799, 0.1651, 0.1527, 0.1419, 0.1326, 0.1244, 1.2490,
0.9828, 0.7854, 0.6435, 0.5404, 0.4636, 0.4049, 0.3588, 0.3218, 0.2915, 0.2663, 0.2450, 0.2268, 0.2111, 0.1974, 0.1854, 1.3258,
1.1072, 0.9273, 0.7854, 0.6747, 0.5880, 0.5191, 0.4636, 0.4182, 0.3805, 0.3488, 0.3218, 0.2985, 0.2783, 0.2606, 0.2450, 1.3734,
1.1903, 1.0304, 0.8961, 0.7854, 0.6947, 0.6203, 0.5586, 0.5071, 0.4636, 0.4266, 0.3948, 0.3672, 0.3430, 0.3218, 0.3029, 1.4057,
1.2490, 1.1072, 0.9828, 0.8761, 0.7854, 0.7086, 0.6435, 0.5880, 0.5404, 0.4993, 0.4636, 0.4324, 0.4049, 0.3805, 0.3588, 1.4289,
1.2925, 1.1659, 1.0517, 0.9505, 0.8622, 0.7854, 0.7188, 0.6610, 0.6107, 0.5667, 0.5281, 0.4939, 0.4636, 0.4366, 0.4124, 1.4464,
1.3258, 1.2120, 1.1072, 1.0122, 0.9273, 0.8520, 0.7854, 0.7267, 0.6747, 0.6288, 0.5880, 0.5517, 0.5191, 0.4899, 0.4636, 1.4601,
1.3521, 1.2490, 1.1526, 1.0637, 0.9828, 0.9098, 0.8441, 0.7854, 0.7328, 0.6857, 0.6435, 0.6055, 0.5713, 0.5404, 0.5124, 1.4711,
1.3734, 1.2793, 1.1903, 1.1072, 1.0304, 0.9601, 0.8961, 0.8380, 0.7854, 0.7378, 0.6947, 0.6557, 0.6203, 0.5880, 0.5586, 1.4801,
1.3909, 1.3045, 1.2220, 1.1442, 1.0715, 1.0041, 0.9420, 0.8851, 0.8330, 0.7854, 0.7419, 0.7023, 0.6660, 0.6328, 0.6023, 1.4877,
1.4057, 1.3258, 1.2490, 1.1760, 1.1072, 1.0427, 0.9828, 0.9273, 0.8761, 0.8289, 0.7854, 0.7454, 0.7086, 0.6747, 0.6435, 1.4940,
1.4182, 1.3440, 1.2723, 1.2036, 1.1384, 1.0769, 1.0191, 0.9653, 0.9151, 0.8685, 0.8254, 0.7854, 0.7484, 0.7141, 0.6823, 1.4995,
1.4289, 1.3597, 1.2925, 1.2278, 1.1659, 1.1072, 1.0517, 0.9995, 0.9505, 0.9048, 0.8622, 0.8224, 0.7854, 0.7509, 0.7188, 1.5042,
1.4382, 1.3734, 1.3102, 1.2490, 1.1903, 1.1342, 1.0809, 1.0304, 0.9828, 0.9380, 0.8961, 0.8567, 0.8199, 0.7854, 0.7531, 1.5084,
1.4464, 1.3854, 1.3258, 1.2679, 1.2120, 1.1584, 1.1072, 1.0584, 1.0122, 0.9685, 0.9273, 0.8885, 0.8520, 0.8177, 0.7854);

Begin
	process (clk, enable, dx, dy)
    begin
        if rising_edge(clk) then
            if enable = '1' then
                magnit <= mem((integer(dx)-1) * 16 + integer(dy)-1);
                angle  <= mem(256 + (integer(dx)-1) * 16 + integer(dy)-1);
            end if;
        end if;
    end process;
End Behavioral;

